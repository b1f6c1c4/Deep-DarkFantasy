module top(
   input clk_i_p,
   input clk_i_n,
   output [3:0] led_o,
   input [3:0] button_ni,

   // HDMI in
   inout vout_scl_io,
   inout vout_sda_io,
   output vout_clk_o,
   output reg vout_de_o,
   output reg vout_hs_o,
   output reg vout_vs_o,
   output reg [23:0] vout_data_o,

   // HDMI out
   inout vin_scl_io,
   inout vin_sda_io,
   input vin_clk_i,
   output vin_rst_no,
   input vin_de_i,
   input vin_hs_i,
   input vin_vs_i,
   input [23:0] vin_data_i,

   output fan_no
);

   localparam WN = 1920;
   localparam KN = 10;
   localparam DELAYS = WN*KN+1;

   wire rst_n = button_ni[0];

   assign fan_no = 0;

   wire clk_video; // 148.571MHz
   wire clk_i2c; // 100MHz
   wire pll_locked;
   sys_pll i_sys_pll (
      .clk_in1_p (clk_i_p),
      .clk_in1_n (clk_i_n),
      .reset (~rst_n),
      .clk_out1 (clk_video),
      .clk_out2 (clk_i2c),
      .locked (pll_locked)
   );

   // HDMI in
   assign vin_rst_no = rst_n;
   sil9013 i_sil9013 (
      .clk_i (clk_i2c),
      .rst_ni (rst_n),
      .vin_scl_io,
      .vin_sda_io
   );
   reg vin_hs, vin_vs, vin_de;
   reg [23:0] vin_data;
   always @(posedge vin_clk_i) begin
      vin_hs <= vin_hs_i;
      vin_vs <= vin_vs_i;
      vin_de <= vin_de_i;
      vin_data <= vin_data_i;
   end

   // Gray calculation
   wire [7:0] gray;
   rgb_to_gray i_rgb_to_gray (
      .r_i(vin_data[23:16]),
      .g_i(vin_data[15:8]),
      .b_i(vin_data[7:0]),
      .k_o(gray)
   );

   // Block buffer
   reg vin_hs_r;
   reg [31:0] h_cur, hb_cur, vp_cur;
   always @(posedge vin_clk_i) begin
      if (vin_vs) begin
         h_cur <= 0;
         hb_cur <= 0;
         vp_cur <= 0;
         vin_hs_r <= 0;
      end else begin
         vin_hs_r <= vin_hs;
         if (vin_hs && ~vin_hs_r) begin
            vp_cur <= (vp_cur == KN-1) ? 0 : vp_cur + 1;
         end
         if (vin_de) begin
            if (h_cur == KN-1) begin
               h_cur <= 0;
               hb_cur <= hb_cur + 1;
            end else begin
               h_cur <= h_cur + 1;
            end
         end
      end
   end

   reg [31:0] blk_buf_a[0:WN/KN-1];
   reg [31:0] blk_buf_b[0:WN/KN-1];
   genvar i;
   generate
      for (i = 0; i < WN/KN; i = i + 1) begin : gen_buffer
         always @(posedge vin_clk_i) begin
            if (vin_vs) begin
               blk_buf_a[i] <= 0;
               blk_buf_b[i] <= 0;
            end else if (vin_hs && ~vin_hs_r && vp_cur == KN-1) begin
               blk_buf_a[i] <= blk_buf_b[i];
               blk_buf_b[i] <= 0;
            end else if (vin_de && i == hb_cur) begin
               blk_buf_b[i] <= blk_buf_b[i] + gray;
            end
         end
      end
   endgenerate

   // Extra stages
   reg [26:0] delay[0:DELAYS-1];
   generate
      for (i = 0; i < DELAYS-1; i = i + 1) begin : gen_delay
         always @(posedge vin_clk_i, negedge rst_n) begin
            if (~rst_n) begin
               delay[i] <= 0;
            end else begin
               delay[i] <= delay[i + 1];
            end
         end
      end
   endgenerate
   always @(posedge vin_clk_i, negedge rst_n) begin
      if (~rst_n) begin
         delay[DELAYS-1] <= 0;
      end else begin
         delay[DELAYS-1] <= {vin_hs, vin_vs, vin_de, vin_data};
      end
   end

   // Output selection
   wire [31:0] active_blk = blk_buf_a[hb_cur];
   wire active_light = active_blk > (KN * KN * 255 / 2);
   assign vout_clk_o = vin_clk_i;
   reg vout_hs;
   reg vout_vs;
   reg vout_de;
   reg [23:0] vout_data;
   always @(*) begin
      if (button_ni[1]) begin
         vout_hs = delay[0][26];
         vout_vs = delay[0][25];
         vout_de = delay[0][24];
         vout_data = {24{active_light}} ^ delay[0][23:0];
      end else begin
         vout_hs = vin_hs;
         vout_vs = vin_hs;
         vout_de = vin_de;
         vout_data = vin_data;
      end
   end

   // HDMI out
   adv7511 i_adv7511 (
      .clk_i (clk_i2c),
      .rst_ni (rst_n),
      .vout_scl_io,
      .vout_sda_io
   );
   always @(posedge vin_clk_i) begin
      vout_hs_o <= vout_hs;
      vout_vs_o <= vout_vs;
      vout_de_o <= vout_de;
      vout_data_o <= vout_data;
   end

endmodule
