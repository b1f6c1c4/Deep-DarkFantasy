module rgb_to_gray (
   input [7:0] r_i,
   input [7:0] g_i,
   input [7:0] b_i,
   output reg [7:0] k_o
);

   reg [21:0] Y;
   always @(*) begin
      Y = 0;
      Y = Y + 2126 * {1'b0,r_i};
      Y = Y + 7152 * {1'b0,g_i};
      Y = Y + 0722 * {1'b0,b_i};
   end

   always @(*) begin
      case (Y[21:12])
         10'd0: k_o = 8'd0;
         10'd1: k_o = 8'd0;
         10'd2: k_o = 8'd1;
         10'd3: k_o = 8'd1;
         10'd4: k_o = 8'd2;
         10'd5: k_o = 8'd2;
         10'd6: k_o = 8'd2;
         10'd7: k_o = 8'd3;
         10'd8: k_o = 8'd3;
         10'd9: k_o = 8'd4;
         10'd10: k_o = 8'd4;
         10'd11: k_o = 8'd5;
         10'd12: k_o = 8'd5;
         10'd13: k_o = 8'd5;
         10'd14: k_o = 8'd6;
         10'd15: k_o = 8'd6;
         10'd16: k_o = 8'd7;
         10'd17: k_o = 8'd7;
         10'd18: k_o = 8'd7;
         10'd19: k_o = 8'd8;
         10'd20: k_o = 8'd8;
         10'd21: k_o = 8'd9;
         10'd22: k_o = 8'd9;
         10'd23: k_o = 8'd9;
         10'd24: k_o = 8'd10;
         10'd25: k_o = 8'd10;
         10'd26: k_o = 8'd11;
         10'd27: k_o = 8'd11;
         10'd28: k_o = 8'd11;
         10'd29: k_o = 8'd12;
         10'd30: k_o = 8'd12;
         10'd31: k_o = 8'd13;
         10'd32: k_o = 8'd13;
         10'd33: k_o = 8'd14;
         10'd34: k_o = 8'd14;
         10'd35: k_o = 8'd14;
         10'd36: k_o = 8'd15;
         10'd37: k_o = 8'd15;
         10'd38: k_o = 8'd16;
         10'd39: k_o = 8'd16;
         10'd40: k_o = 8'd16;
         10'd41: k_o = 8'd17;
         10'd42: k_o = 8'd17;
         10'd43: k_o = 8'd18;
         10'd44: k_o = 8'd18;
         10'd45: k_o = 8'd18;
         10'd46: k_o = 8'd19;
         10'd47: k_o = 8'd19;
         10'd48: k_o = 8'd20;
         10'd49: k_o = 8'd20;
         10'd50: k_o = 8'd20;
         10'd51: k_o = 8'd21;
         10'd52: k_o = 8'd21;
         10'd53: k_o = 8'd22;
         10'd54: k_o = 8'd22;
         10'd55: k_o = 8'd23;
         10'd56: k_o = 8'd23;
         10'd57: k_o = 8'd23;
         10'd58: k_o = 8'd24;
         10'd59: k_o = 8'd24;
         10'd60: k_o = 8'd25;
         10'd61: k_o = 8'd25;
         10'd62: k_o = 8'd25;
         10'd63: k_o = 8'd26;
         10'd64: k_o = 8'd26;
         10'd65: k_o = 8'd27;
         10'd66: k_o = 8'd27;
         10'd67: k_o = 8'd27;
         10'd68: k_o = 8'd28;
         10'd69: k_o = 8'd28;
         10'd70: k_o = 8'd29;
         10'd71: k_o = 8'd29;
         10'd72: k_o = 8'd29;
         10'd73: k_o = 8'd30;
         10'd74: k_o = 8'd30;
         10'd75: k_o = 8'd31;
         10'd76: k_o = 8'd31;
         10'd77: k_o = 8'd32;
         10'd78: k_o = 8'd32;
         10'd79: k_o = 8'd32;
         10'd80: k_o = 8'd33;
         10'd81: k_o = 8'd33;
         10'd82: k_o = 8'd34;
         10'd83: k_o = 8'd34;
         10'd84: k_o = 8'd34;
         10'd85: k_o = 8'd35;
         10'd86: k_o = 8'd35;
         10'd87: k_o = 8'd36;
         10'd88: k_o = 8'd36;
         10'd89: k_o = 8'd36;
         10'd90: k_o = 8'd37;
         10'd91: k_o = 8'd37;
         10'd92: k_o = 8'd38;
         10'd93: k_o = 8'd38;
         10'd94: k_o = 8'd39;
         10'd95: k_o = 8'd39;
         10'd96: k_o = 8'd39;
         10'd97: k_o = 8'd40;
         10'd98: k_o = 8'd40;
         10'd99: k_o = 8'd41;
         10'd100: k_o = 8'd41;
         10'd101: k_o = 8'd41;
         10'd102: k_o = 8'd42;
         10'd103: k_o = 8'd42;
         10'd104: k_o = 8'd43;
         10'd105: k_o = 8'd43;
         10'd106: k_o = 8'd43;
         10'd107: k_o = 8'd44;
         10'd108: k_o = 8'd44;
         10'd109: k_o = 8'd45;
         10'd110: k_o = 8'd45;
         10'd111: k_o = 8'd45;
         10'd112: k_o = 8'd46;
         10'd113: k_o = 8'd46;
         10'd114: k_o = 8'd47;
         10'd115: k_o = 8'd47;
         10'd116: k_o = 8'd48;
         10'd117: k_o = 8'd48;
         10'd118: k_o = 8'd48;
         10'd119: k_o = 8'd49;
         10'd120: k_o = 8'd49;
         10'd121: k_o = 8'd50;
         10'd122: k_o = 8'd50;
         10'd123: k_o = 8'd50;
         10'd124: k_o = 8'd51;
         10'd125: k_o = 8'd51;
         10'd126: k_o = 8'd52;
         10'd127: k_o = 8'd52;
         10'd128: k_o = 8'd52;
         10'd129: k_o = 8'd53;
         10'd130: k_o = 8'd53;
         10'd131: k_o = 8'd54;
         10'd132: k_o = 8'd54;
         10'd133: k_o = 8'd54;
         10'd134: k_o = 8'd55;
         10'd135: k_o = 8'd55;
         10'd136: k_o = 8'd56;
         10'd137: k_o = 8'd56;
         10'd138: k_o = 8'd57;
         10'd139: k_o = 8'd57;
         10'd140: k_o = 8'd57;
         10'd141: k_o = 8'd58;
         10'd142: k_o = 8'd58;
         10'd143: k_o = 8'd59;
         10'd144: k_o = 8'd59;
         10'd145: k_o = 8'd59;
         10'd146: k_o = 8'd60;
         10'd147: k_o = 8'd60;
         10'd148: k_o = 8'd61;
         10'd149: k_o = 8'd61;
         10'd150: k_o = 8'd61;
         10'd151: k_o = 8'd62;
         10'd152: k_o = 8'd62;
         10'd153: k_o = 8'd63;
         10'd154: k_o = 8'd63;
         10'd155: k_o = 8'd63;
         10'd156: k_o = 8'd64;
         10'd157: k_o = 8'd64;
         10'd158: k_o = 8'd65;
         10'd159: k_o = 8'd65;
         10'd160: k_o = 8'd66;
         10'd161: k_o = 8'd66;
         10'd162: k_o = 8'd66;
         10'd163: k_o = 8'd67;
         10'd164: k_o = 8'd67;
         10'd165: k_o = 8'd68;
         10'd166: k_o = 8'd68;
         10'd167: k_o = 8'd68;
         10'd168: k_o = 8'd69;
         10'd169: k_o = 8'd69;
         10'd170: k_o = 8'd70;
         10'd171: k_o = 8'd70;
         10'd172: k_o = 8'd70;
         10'd173: k_o = 8'd71;
         10'd174: k_o = 8'd71;
         10'd175: k_o = 8'd72;
         10'd176: k_o = 8'd72;
         10'd177: k_o = 8'd72;
         10'd178: k_o = 8'd73;
         10'd179: k_o = 8'd73;
         10'd180: k_o = 8'd74;
         10'd181: k_o = 8'd74;
         10'd182: k_o = 8'd75;
         10'd183: k_o = 8'd75;
         10'd184: k_o = 8'd75;
         10'd185: k_o = 8'd76;
         10'd186: k_o = 8'd76;
         10'd187: k_o = 8'd77;
         10'd188: k_o = 8'd77;
         10'd189: k_o = 8'd77;
         10'd190: k_o = 8'd78;
         10'd191: k_o = 8'd78;
         10'd192: k_o = 8'd79;
         10'd193: k_o = 8'd79;
         10'd194: k_o = 8'd79;
         10'd195: k_o = 8'd80;
         10'd196: k_o = 8'd80;
         10'd197: k_o = 8'd81;
         10'd198: k_o = 8'd81;
         10'd199: k_o = 8'd82;
         10'd200: k_o = 8'd82;
         10'd201: k_o = 8'd82;
         10'd202: k_o = 8'd83;
         10'd203: k_o = 8'd83;
         10'd204: k_o = 8'd84;
         10'd205: k_o = 8'd84;
         10'd206: k_o = 8'd84;
         10'd207: k_o = 8'd85;
         10'd208: k_o = 8'd85;
         10'd209: k_o = 8'd86;
         10'd210: k_o = 8'd86;
         10'd211: k_o = 8'd86;
         10'd212: k_o = 8'd87;
         10'd213: k_o = 8'd87;
         10'd214: k_o = 8'd88;
         10'd215: k_o = 8'd88;
         10'd216: k_o = 8'd88;
         10'd217: k_o = 8'd89;
         10'd218: k_o = 8'd89;
         10'd219: k_o = 8'd90;
         10'd220: k_o = 8'd90;
         10'd221: k_o = 8'd91;
         10'd222: k_o = 8'd91;
         10'd223: k_o = 8'd91;
         10'd224: k_o = 8'd92;
         10'd225: k_o = 8'd92;
         10'd226: k_o = 8'd93;
         10'd227: k_o = 8'd93;
         10'd228: k_o = 8'd93;
         10'd229: k_o = 8'd94;
         10'd230: k_o = 8'd94;
         10'd231: k_o = 8'd95;
         10'd232: k_o = 8'd95;
         10'd233: k_o = 8'd95;
         10'd234: k_o = 8'd96;
         10'd235: k_o = 8'd96;
         10'd236: k_o = 8'd97;
         10'd237: k_o = 8'd97;
         10'd238: k_o = 8'd97;
         10'd239: k_o = 8'd98;
         10'd240: k_o = 8'd98;
         10'd241: k_o = 8'd99;
         10'd242: k_o = 8'd99;
         10'd243: k_o = 8'd100;
         10'd244: k_o = 8'd100;
         10'd245: k_o = 8'd100;
         10'd246: k_o = 8'd101;
         10'd247: k_o = 8'd101;
         10'd248: k_o = 8'd102;
         10'd249: k_o = 8'd102;
         10'd250: k_o = 8'd102;
         10'd251: k_o = 8'd103;
         10'd252: k_o = 8'd103;
         10'd253: k_o = 8'd104;
         10'd254: k_o = 8'd104;
         10'd255: k_o = 8'd104;
         10'd256: k_o = 8'd105;
         10'd257: k_o = 8'd105;
         10'd258: k_o = 8'd106;
         10'd259: k_o = 8'd106;
         10'd260: k_o = 8'd106;
         10'd261: k_o = 8'd107;
         10'd262: k_o = 8'd107;
         10'd263: k_o = 8'd108;
         10'd264: k_o = 8'd108;
         10'd265: k_o = 8'd109;
         10'd266: k_o = 8'd109;
         10'd267: k_o = 8'd109;
         10'd268: k_o = 8'd110;
         10'd269: k_o = 8'd110;
         10'd270: k_o = 8'd111;
         10'd271: k_o = 8'd111;
         10'd272: k_o = 8'd111;
         10'd273: k_o = 8'd112;
         10'd274: k_o = 8'd112;
         10'd275: k_o = 8'd113;
         10'd276: k_o = 8'd113;
         10'd277: k_o = 8'd113;
         10'd278: k_o = 8'd114;
         10'd279: k_o = 8'd114;
         10'd280: k_o = 8'd115;
         10'd281: k_o = 8'd115;
         10'd282: k_o = 8'd116;
         10'd283: k_o = 8'd116;
         10'd284: k_o = 8'd116;
         10'd285: k_o = 8'd117;
         10'd286: k_o = 8'd117;
         10'd287: k_o = 8'd118;
         10'd288: k_o = 8'd118;
         10'd289: k_o = 8'd118;
         10'd290: k_o = 8'd119;
         10'd291: k_o = 8'd119;
         10'd292: k_o = 8'd120;
         10'd293: k_o = 8'd120;
         10'd294: k_o = 8'd120;
         10'd295: k_o = 8'd121;
         10'd296: k_o = 8'd121;
         10'd297: k_o = 8'd122;
         10'd298: k_o = 8'd122;
         10'd299: k_o = 8'd122;
         10'd300: k_o = 8'd123;
         10'd301: k_o = 8'd123;
         10'd302: k_o = 8'd124;
         10'd303: k_o = 8'd124;
         10'd304: k_o = 8'd125;
         10'd305: k_o = 8'd125;
         10'd306: k_o = 8'd125;
         10'd307: k_o = 8'd126;
         10'd308: k_o = 8'd126;
         10'd309: k_o = 8'd127;
         10'd310: k_o = 8'd127;
         10'd311: k_o = 8'd127;
         10'd312: k_o = 8'd128;
         10'd313: k_o = 8'd128;
         10'd314: k_o = 8'd129;
         10'd315: k_o = 8'd129;
         10'd316: k_o = 8'd129;
         10'd317: k_o = 8'd130;
         10'd318: k_o = 8'd130;
         10'd319: k_o = 8'd131;
         10'd320: k_o = 8'd131;
         10'd321: k_o = 8'd131;
         10'd322: k_o = 8'd132;
         10'd323: k_o = 8'd132;
         10'd324: k_o = 8'd133;
         10'd325: k_o = 8'd133;
         10'd326: k_o = 8'd134;
         10'd327: k_o = 8'd134;
         10'd328: k_o = 8'd134;
         10'd329: k_o = 8'd135;
         10'd330: k_o = 8'd135;
         10'd331: k_o = 8'd136;
         10'd332: k_o = 8'd136;
         10'd333: k_o = 8'd136;
         10'd334: k_o = 8'd137;
         10'd335: k_o = 8'd137;
         10'd336: k_o = 8'd138;
         10'd337: k_o = 8'd138;
         10'd338: k_o = 8'd138;
         10'd339: k_o = 8'd139;
         10'd340: k_o = 8'd139;
         10'd341: k_o = 8'd140;
         10'd342: k_o = 8'd140;
         10'd343: k_o = 8'd140;
         10'd344: k_o = 8'd141;
         10'd345: k_o = 8'd141;
         10'd346: k_o = 8'd142;
         10'd347: k_o = 8'd142;
         10'd348: k_o = 8'd143;
         10'd349: k_o = 8'd143;
         10'd350: k_o = 8'd143;
         10'd351: k_o = 8'd144;
         10'd352: k_o = 8'd144;
         10'd353: k_o = 8'd145;
         10'd354: k_o = 8'd145;
         10'd355: k_o = 8'd145;
         10'd356: k_o = 8'd146;
         10'd357: k_o = 8'd146;
         10'd358: k_o = 8'd147;
         10'd359: k_o = 8'd147;
         10'd360: k_o = 8'd147;
         10'd361: k_o = 8'd148;
         10'd362: k_o = 8'd148;
         10'd363: k_o = 8'd149;
         10'd364: k_o = 8'd149;
         10'd365: k_o = 8'd150;
         10'd366: k_o = 8'd150;
         10'd367: k_o = 8'd150;
         10'd368: k_o = 8'd151;
         10'd369: k_o = 8'd151;
         10'd370: k_o = 8'd152;
         10'd371: k_o = 8'd152;
         10'd372: k_o = 8'd152;
         10'd373: k_o = 8'd153;
         10'd374: k_o = 8'd153;
         10'd375: k_o = 8'd154;
         10'd376: k_o = 8'd154;
         10'd377: k_o = 8'd154;
         10'd378: k_o = 8'd155;
         10'd379: k_o = 8'd155;
         10'd380: k_o = 8'd156;
         10'd381: k_o = 8'd156;
         10'd382: k_o = 8'd156;
         10'd383: k_o = 8'd157;
         10'd384: k_o = 8'd157;
         10'd385: k_o = 8'd158;
         10'd386: k_o = 8'd158;
         10'd387: k_o = 8'd159;
         10'd388: k_o = 8'd159;
         10'd389: k_o = 8'd159;
         10'd390: k_o = 8'd160;
         10'd391: k_o = 8'd160;
         10'd392: k_o = 8'd161;
         10'd393: k_o = 8'd161;
         10'd394: k_o = 8'd161;
         10'd395: k_o = 8'd162;
         10'd396: k_o = 8'd162;
         10'd397: k_o = 8'd163;
         10'd398: k_o = 8'd163;
         10'd399: k_o = 8'd163;
         10'd400: k_o = 8'd164;
         10'd401: k_o = 8'd164;
         10'd402: k_o = 8'd165;
         10'd403: k_o = 8'd165;
         10'd404: k_o = 8'd165;
         10'd405: k_o = 8'd166;
         10'd406: k_o = 8'd166;
         10'd407: k_o = 8'd167;
         10'd408: k_o = 8'd167;
         10'd409: k_o = 8'd168;
         10'd410: k_o = 8'd168;
         10'd411: k_o = 8'd168;
         10'd412: k_o = 8'd169;
         10'd413: k_o = 8'd169;
         10'd414: k_o = 8'd170;
         10'd415: k_o = 8'd170;
         10'd416: k_o = 8'd170;
         10'd417: k_o = 8'd171;
         10'd418: k_o = 8'd171;
         10'd419: k_o = 8'd172;
         10'd420: k_o = 8'd172;
         10'd421: k_o = 8'd172;
         10'd422: k_o = 8'd173;
         10'd423: k_o = 8'd173;
         10'd424: k_o = 8'd174;
         10'd425: k_o = 8'd174;
         10'd426: k_o = 8'd174;
         10'd427: k_o = 8'd175;
         10'd428: k_o = 8'd175;
         10'd429: k_o = 8'd176;
         10'd430: k_o = 8'd176;
         10'd431: k_o = 8'd177;
         10'd432: k_o = 8'd177;
         10'd433: k_o = 8'd177;
         10'd434: k_o = 8'd178;
         10'd435: k_o = 8'd178;
         10'd436: k_o = 8'd179;
         10'd437: k_o = 8'd179;
         10'd438: k_o = 8'd179;
         10'd439: k_o = 8'd180;
         10'd440: k_o = 8'd180;
         10'd441: k_o = 8'd181;
         10'd442: k_o = 8'd181;
         10'd443: k_o = 8'd181;
         10'd444: k_o = 8'd182;
         10'd445: k_o = 8'd182;
         10'd446: k_o = 8'd183;
         10'd447: k_o = 8'd183;
         10'd448: k_o = 8'd184;
         10'd449: k_o = 8'd184;
         10'd450: k_o = 8'd184;
         10'd451: k_o = 8'd185;
         10'd452: k_o = 8'd185;
         10'd453: k_o = 8'd186;
         10'd454: k_o = 8'd186;
         10'd455: k_o = 8'd186;
         10'd456: k_o = 8'd187;
         10'd457: k_o = 8'd187;
         10'd458: k_o = 8'd188;
         10'd459: k_o = 8'd188;
         10'd460: k_o = 8'd188;
         10'd461: k_o = 8'd189;
         10'd462: k_o = 8'd189;
         10'd463: k_o = 8'd190;
         10'd464: k_o = 8'd190;
         10'd465: k_o = 8'd190;
         10'd466: k_o = 8'd191;
         10'd467: k_o = 8'd191;
         10'd468: k_o = 8'd192;
         10'd469: k_o = 8'd192;
         10'd470: k_o = 8'd193;
         10'd471: k_o = 8'd193;
         10'd472: k_o = 8'd193;
         10'd473: k_o = 8'd194;
         10'd474: k_o = 8'd194;
         10'd475: k_o = 8'd195;
         10'd476: k_o = 8'd195;
         10'd477: k_o = 8'd195;
         10'd478: k_o = 8'd196;
         10'd479: k_o = 8'd196;
         10'd480: k_o = 8'd197;
         10'd481: k_o = 8'd197;
         10'd482: k_o = 8'd197;
         10'd483: k_o = 8'd198;
         10'd484: k_o = 8'd198;
         10'd485: k_o = 8'd199;
         10'd486: k_o = 8'd199;
         10'd487: k_o = 8'd199;
         10'd488: k_o = 8'd200;
         10'd489: k_o = 8'd200;
         10'd490: k_o = 8'd201;
         10'd491: k_o = 8'd201;
         10'd492: k_o = 8'd202;
         10'd493: k_o = 8'd202;
         10'd494: k_o = 8'd202;
         10'd495: k_o = 8'd203;
         10'd496: k_o = 8'd203;
         10'd497: k_o = 8'd204;
         10'd498: k_o = 8'd204;
         10'd499: k_o = 8'd204;
         10'd500: k_o = 8'd205;
         10'd501: k_o = 8'd205;
         10'd502: k_o = 8'd206;
         10'd503: k_o = 8'd206;
         10'd504: k_o = 8'd206;
         10'd505: k_o = 8'd207;
         10'd506: k_o = 8'd207;
         10'd507: k_o = 8'd208;
         10'd508: k_o = 8'd208;
         10'd509: k_o = 8'd208;
         10'd510: k_o = 8'd209;
         10'd511: k_o = 8'd209;
         10'd512: k_o = 8'd210;
         10'd513: k_o = 8'd210;
         10'd514: k_o = 8'd211;
         10'd515: k_o = 8'd211;
         10'd516: k_o = 8'd211;
         10'd517: k_o = 8'd212;
         10'd518: k_o = 8'd212;
         10'd519: k_o = 8'd213;
         10'd520: k_o = 8'd213;
         10'd521: k_o = 8'd213;
         10'd522: k_o = 8'd214;
         10'd523: k_o = 8'd214;
         10'd524: k_o = 8'd215;
         10'd525: k_o = 8'd215;
         10'd526: k_o = 8'd215;
         10'd527: k_o = 8'd216;
         10'd528: k_o = 8'd216;
         10'd529: k_o = 8'd217;
         10'd530: k_o = 8'd217;
         10'd531: k_o = 8'd217;
         10'd532: k_o = 8'd218;
         10'd533: k_o = 8'd218;
         10'd534: k_o = 8'd219;
         10'd535: k_o = 8'd219;
         10'd536: k_o = 8'd220;
         10'd537: k_o = 8'd220;
         10'd538: k_o = 8'd220;
         10'd539: k_o = 8'd221;
         10'd540: k_o = 8'd221;
         10'd541: k_o = 8'd222;
         10'd542: k_o = 8'd222;
         10'd543: k_o = 8'd222;
         10'd544: k_o = 8'd223;
         10'd545: k_o = 8'd223;
         10'd546: k_o = 8'd224;
         10'd547: k_o = 8'd224;
         10'd548: k_o = 8'd224;
         10'd549: k_o = 8'd225;
         10'd550: k_o = 8'd225;
         10'd551: k_o = 8'd226;
         10'd552: k_o = 8'd226;
         10'd553: k_o = 8'd227;
         10'd554: k_o = 8'd227;
         10'd555: k_o = 8'd227;
         10'd556: k_o = 8'd228;
         10'd557: k_o = 8'd228;
         10'd558: k_o = 8'd229;
         10'd559: k_o = 8'd229;
         10'd560: k_o = 8'd229;
         10'd561: k_o = 8'd230;
         10'd562: k_o = 8'd230;
         10'd563: k_o = 8'd231;
         10'd564: k_o = 8'd231;
         10'd565: k_o = 8'd231;
         10'd566: k_o = 8'd232;
         10'd567: k_o = 8'd232;
         10'd568: k_o = 8'd233;
         10'd569: k_o = 8'd233;
         10'd570: k_o = 8'd233;
         10'd571: k_o = 8'd234;
         10'd572: k_o = 8'd234;
         10'd573: k_o = 8'd235;
         10'd574: k_o = 8'd235;
         10'd575: k_o = 8'd236;
         10'd576: k_o = 8'd236;
         10'd577: k_o = 8'd236;
         10'd578: k_o = 8'd237;
         10'd579: k_o = 8'd237;
         10'd580: k_o = 8'd238;
         10'd581: k_o = 8'd238;
         10'd582: k_o = 8'd238;
         10'd583: k_o = 8'd239;
         10'd584: k_o = 8'd239;
         10'd585: k_o = 8'd240;
         10'd586: k_o = 8'd240;
         10'd587: k_o = 8'd240;
         10'd588: k_o = 8'd241;
         10'd589: k_o = 8'd241;
         10'd590: k_o = 8'd242;
         10'd591: k_o = 8'd242;
         10'd592: k_o = 8'd242;
         10'd593: k_o = 8'd243;
         10'd594: k_o = 8'd243;
         10'd595: k_o = 8'd244;
         10'd596: k_o = 8'd244;
         10'd597: k_o = 8'd245;
         10'd598: k_o = 8'd245;
         10'd599: k_o = 8'd245;
         10'd600: k_o = 8'd246;
         10'd601: k_o = 8'd246;
         10'd602: k_o = 8'd247;
         10'd603: k_o = 8'd247;
         10'd604: k_o = 8'd247;
         10'd605: k_o = 8'd248;
         10'd606: k_o = 8'd248;
         10'd607: k_o = 8'd249;
         10'd608: k_o = 8'd249;
         10'd609: k_o = 8'd249;
         10'd610: k_o = 8'd250;
         10'd611: k_o = 8'd250;
         10'd612: k_o = 8'd251;
         10'd613: k_o = 8'd251;
         10'd614: k_o = 8'd251;
         10'd615: k_o = 8'd252;
         10'd616: k_o = 8'd252;
         10'd617: k_o = 8'd253;
         10'd618: k_o = 8'd253;
         10'd619: k_o = 8'd254;
         10'd620: k_o = 8'd254;
         10'd621: k_o = 8'd254;
         default: k_o = 8'd255;
      endcase
   end

endmodule
