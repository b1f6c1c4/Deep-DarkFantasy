module mem (
   input clk_i_p,
   input clk_i_n,
   input rst_ni,
   input step_i,
   input [23:0] data_i,
   output [23:0] data_o
);

   // TODO

endmodule
